// Copyright 2025 Maktab-e-Digital Systems Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description:
// This module implements address matching for NAPOT mode.
//
// Inputs:
// - addr       : [31:0] (unsigned) Base address of the memory region to be accessed.
// - addr_n     : [31:0] (unsigned) Value of the nth PMP address register.
// - size       : [1:0]             Size of the memory access (00: byte, 01: half-word, 11: word).
//
// Output:
// - napot_out  : [0:0]             High if the memory region is supposedly protected by the Nth PMP entry; low otherwise.
//
// Dependencies:
// There are no dependancies. 
//
// Author: Muhammad Boota, Muhammad Furrukh
// Date:

module napot (
    input logic unsigned [31:0] addr, addr_n,
    input logic          [1:0]  size,
    output logic                napot_out
);

logic [5:0]  position;
logic [31:0] ones, base,offset;

assign ones   = (~(32'b0) << position + 1);
assign base   = (addr_n & (ones));
assign offset = (32'h8<<position);
always_comb begin
    napot_out = (( (addr + size) <= (base + offset - 1) ) && ( base <= addr ));
end



always_comb begin :priority_circuit
    casez (addr_n)  // casez allows ? for don't-care bits
        32'b???????????????????????????????0: position = 6'd0;
        32'b??????????????????????????????01: position = 6'd1;
        32'b?????????????????????????????011: position = 6'd2;
        32'b????????????????????????????0111: position = 6'd3;
        32'b???????????????????????????01111: position = 6'd4;
        32'b??????????????????????????011111: position = 6'd5;
        32'b?????????????????????????0111111: position = 6'd6;
        32'b????????????????????????01111111: position = 6'd7;
        32'b???????????????????????011111111: position = 6'd8;
        32'b??????????????????????0111111111: position = 6'd9;
        32'b?????????????????????01111111111: position = 6'd10;
        32'b????????????????????011111111111: position = 6'd11;
        32'b???????????????????0111111111111: position = 6'd12;
        32'b??????????????????01111111111111: position = 6'd13;
        32'b?????????????????011111111111111: position = 6'd14;
        32'b????????????????0111111111111111: position = 6'd15;
        32'b???????????????01111111111111111: position = 6'd16;
        32'b??????????????011111111111111111: position = 6'd17;
        32'b?????????????0111111111111111111: position = 6'd18;
        32'b????????????01111111111111111111: position = 6'd19;
        32'b???????????011111111111111111111: position = 6'd20;
        32'b??????????0111111111111111111111: position = 6'd21;
        32'b?????????01111111111111111111111: position = 6'd22;
        32'b????????011111111111111111111111: position = 6'd23;
        32'b???????0111111111111111111111111: position = 6'd24;
        32'b??????01111111111111111111111111: position = 6'd25;
        32'b?????011111111111111111111111111: position = 6'd26;
        32'b????0111111111111111111111111111: position = 6'd27;
        32'b???01111111111111111111111111111: position = 6'd28;
        32'b??011111111111111111111111111111: position = 6'd29;
        32'b?0111111111111111111111111111111: position = 6'd30;
        32'b01111111111111111111111111111111: position = 6'd31;
        32'b11111111111111111111111111111111: position = 6'd32;
        default:                              position = 6'd0;  // When no bits are set
    endcase
end
endmodule